//Verilog HDL code for pre midterm Problem 12
//Made by: Jhury Kevin P. Lastre
//Date: 9/28/2022

module Problem12 (W, X, Y, Z, D);

	input W, X, Y, Z;
	output D;
	
	wire s1, s2, s3, s4, s5, s6, s7;
	
	not G1 (s1, Z);
	or  G2 (s2, s1, Y);
	not G3 (s3, X);
	and G4 (s4, W, s3);
	not G5 (s5, W);
	and G6 (s6, X, s5);
	or  G7 (s7, s4, s6);
	and G8 (D, s7, s2);

endmodule